module ControlUnit (opcode,func,aluop,regdst,memtoreg,alusrc,regwrite,memread,memwrite,branch,jump,pcsrc);
    input [5:0] opcode,func;
    output reg [2:0] aluop;
    output reg [1:0] regdst,memtoreg;
    output reg alusrc,regwrite,memread,memwrite,branch,jump,pcsrc;
    always @(opcode or func) begin
        if(!opcode) begin
            case(func)
                6'b000000 : begin
                    aluop=3'b000;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b000001 : begin
                    aluop=3'b001;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b000010 : begin
                    aluop=3'b010;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b000011 : begin
                    aluop=3'b011;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b000100 : begin
                    aluop=3'b100;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b000101 : begin
                    aluop=3'b101;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b000110 : begin
                    aluop=3'b110;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b000111 :begin
                    aluop=3'b111;
                    alusrc=0;
                    regdst=2'b01;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b001000 :begin
                    regwrite=0;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=1;
                end
            endcase
        end
        else begin
            case(opcode)
                6'b010000:begin
                    aluop=3'b000;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b010001:begin
                    aluop=3'b001;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b010010:begin
                    aluop=3'b010;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b010011:begin
                    aluop=3'b011;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b010100:begin
                    aluop=3'b100;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b010101:begin
                    aluop=3'b101;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b010110:begin
                    aluop=3'b110;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b010111:begin
                    aluop=3'b111;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b00;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b100011:begin
                    aluop=3'b011;
                    alusrc=1;
                    regdst=2'b00;
                    memtoreg=2'b01;
                    regwrite=1;
                    memread=1;
                    memwrite=0;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b101011:begin
                    aluop=3'b011;
                    alusrc=1;
                    regwrite=0;
                    memread=0;
                    memwrite=1;
                    branch=0;
                    jump=0;
                    pcsrc=0;
                end
                6'b110000:begin
                    regwrite=0;
                    memread=0;
                    memwrite=0;
                    branch=1;
                    jump=0;
                    pcsrc=0;
                end
                6'b110001:begin
                    regwrite=0;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=1;
                    pcsrc=1;
                end
                6'b110011:begin
                    regdst=2'b10;
                    memtoreg=2'b10;
                    regwrite=1;
                    memread=0;
                    memwrite=0;
                    branch=0;
                    jump=1;
                    pcsrc=1;
                end
            endcase
        end
    end
endmodule